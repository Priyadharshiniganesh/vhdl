
entity to1 is
  
end entity to1;

architecture sim of to1 is

begin  -- architecture sim

process is
begin  -- process

  report "Hello World";
  wait;
 
  
end process;

end architecture sim;
